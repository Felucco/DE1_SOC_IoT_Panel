module Graph_TH_Handler (
	input [4:0] px_code,
	output [7:0] graph_R, graph_G, graph_B);
	
	s

endmodule